`define rf_fft_impl _hxfcpuabvjh
`define rf_fft_impl_pkg _hxfcpuabvjh_pkg

package _hxfcpuabvjh_pkg;
    parameter BULK_ADDR_WIDTH = 4;
    parameter BULK_BITWIDTH = 256;
    parameter FSM_PER_SLOT = 4;
    parameter INSTR_OPCODE_BITWIDTH = 3;
    parameter IO_ADDR_WIDTH = 16;
    parameter IO_DATA_WIDTH = 256;
    parameter NUM_SLOTS = 16;
    parameter RESOURCE_INSTR_WIDTH = 27;
    parameter RF_DEPTH = 128;
    parameter WORD_ADDR_WIDTH = 7;
    parameter WORD_BITWIDTH = 32;

    typedef struct packed {
        logic _init_addr_sd;
        logic [15:0] _init_addr;
        logic [1:0] _port;
    } dsu_t;

    function static dsu_t unpack_dsu;
        input logic [23:0] instr;
        dsu_t _dsu;
        _dsu._init_addr_sd = instr[23];
        _dsu._init_addr  = instr[22:7];
        _dsu._port  = instr[6:5];
        return _dsu;
    endfunction

    function static logic [23:0] pack_dsu;
        input dsu_t _dsu;
        logic [23:0] instr;

        instr[23] = _dsu._init_addr_sd;
        instr[22:7] = _dsu._init_addr;
        instr[6:5] = _dsu._port;
        return instr;
    endfunction
    typedef struct packed {
        logic [1:0] _port;
        logic [3:0] _level;
        logic [5:0] _iter;
        logic [5:0] _step;
        logic [5:0] _delay;
    } rep_t;

    function static rep_t unpack_rep;
        input logic [23:0] instr;
        rep_t _rep;
        _rep._port  = instr[23:22];
        _rep._level  = instr[21:18];
        _rep._iter  = instr[17:12];
        _rep._step  = instr[11:6];
        _rep._delay  = instr[5:0];
        return _rep;
    endfunction

    function static logic [23:0] pack_rep;
        input rep_t _rep;
        logic [23:0] instr;

        instr[23:22] = _rep._port;
        instr[21:18] = _rep._level;
        instr[17:12] = _rep._iter;
        instr[11:6] = _rep._step;
        instr[5:0] = _rep._delay;
        return instr;
    endfunction
    typedef struct packed {
        logic [1:0] _port;
        logic [11:0] _n_points;
        logic [1:0] _radix;
        logic _n_bu;
        logic _mode;
        logic [5:0] _delay;
    } fft_t;

    function static fft_t unpack_fft;
        input logic [23:0] instr;
        fft_t _fft;
        _fft._port  = instr[23:22];
        _fft._n_points  = instr[21:10];
        _fft._radix  = instr[9:8];
        _fft._n_bu = instr[7];
        _fft._mode = instr[6];
        _fft._delay  = instr[5:0];
        return _fft;
    endfunction

    function static logic [23:0] pack_fft;
        input fft_t _fft;
        logic [23:0] instr;

        instr[23:22] = _fft._port;
        instr[21:10] = _fft._n_points;
        instr[9:8] = _fft._radix;
        instr[7] = _fft._n_bu;
        instr[6] = _fft._mode;
        instr[5:0] = _fft._delay;
        return instr;
    endfunction

    parameter AGU_BITWIDTH = 16;
    parameter DELAY_WIDTH = 5;

endpackage

module _hxfcpuabvjh
import _hxfcpuabvjh_pkg::*;
(
    input  logic clk_0,
    input  logic rst_n_0,
    input  logic instr_en_0,
    input  logic [RESOURCE_INSTR_WIDTH-1:0] instr_0,
    input  logic [3:0] activate_0,
    input  logic [WORD_BITWIDTH-1:0] word_data_in_0,
    output logic [WORD_BITWIDTH-1:0] word_data_out_0,
    input  logic [BULK_BITWIDTH-1:0] bulk_data_in_0,
    output logic [BULK_BITWIDTH-1:0] bulk_data_out_0,
    input  logic clk_1,
    input  logic rst_n_1,
    input  logic instr_en_1,
    input  logic [RESOURCE_INSTR_WIDTH-1:0] instr_1,
    input  logic [3:0] activate_1,
    input  logic [WORD_BITWIDTH-1:0] word_data_in_1,
    output logic [WORD_BITWIDTH-1:0] word_data_out_1,
    input  logic [BULK_BITWIDTH-1:0] bulk_data_in_1,
    output logic [BULK_BITWIDTH-1:0] bulk_data_out_1
);

    logic clk, rst_n;
    assign clk = clk_0;
    assign rst_n = rst_n_0;

    assign bulk_data_out_1 = 0;

    logic [RF_DEPTH-1:0][WORD_BITWIDTH-1:0] memory, memory_next;
    logic bulk_w_en, bulk_r_en;
    logic word_w_en_0, word_r_en_0;
    logic word_w_en_1, word_r_en_1;
    logic [BULK_ADDR_WIDTH-1:0] bulk_w_addr, bulk_r_addr;
    logic [WORD_ADDR_WIDTH-1:0] word_w_addr_0, word_r_addr_0;
    logic [WORD_ADDR_WIDTH-1:0] word_w_addr_1, word_r_addr_1;
    logic [AGU_BITWIDTH-1:0] bulk_w_agu, bulk_r_agu;
    logic [AGU_BITWIDTH-1:0] word_w_agu_0, word_r_agu_0;
    logic [AGU_BITWIDTH-1:0] word_w_agu_1, word_r_agu_1;

    assign bulk_w_addr = bulk_w_agu[BULK_ADDR_WIDTH-1:0];
    assign bulk_r_addr = bulk_r_agu[BULK_ADDR_WIDTH-1:0];
    assign word_w_addr_0 = word_w_agu_0[WORD_ADDR_WIDTH-1:0];
    assign word_r_addr_0 = word_r_agu_0[WORD_ADDR_WIDTH-1:0];
    assign word_w_addr_1 = word_w_agu_1[WORD_ADDR_WIDTH-1:0];
    assign word_r_addr_1 = word_r_agu_1[WORD_ADDR_WIDTH-1:0];

    logic fft_valid;
    logic dsu_valid;
    logic rep_valid;

    logic [DELAY_WIDTH-1:0] delay_0_0, delay_0_1;
    logic [AGU_BITWIDTH-1:0] n_points_0_0, n_points_0_1;
    logic [1:0] radix_0_0, radix_0_1;
    logic n_bu_0_0, n_bu_0_1;
    logic mode_0_0, mode_0_1;

    logic [AGU_BITWIDTH-1:0] step_0_2, step_0_3;
    logic [AGU_BITWIDTH-1:0] delay_0_2, delay_0_3;
    logic [AGU_BITWIDTH-1:0] iter_0_2, iter_0_3;
    logic [AGU_BITWIDTH-1:0] init_addr_0_2, init_addr_0_3;

    logic [DELAY_WIDTH-1:0] delay_1_0, delay_1_1;
    logic [AGU_BITWIDTH-1:0] n_points_1_0, n_points_1_1;
    logic [1:0] radix_1_0, radix_1_1;
    logic n_bu_1_0, n_bu_1_1;
    logic mode_1_0, mode_1_1;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            memory <= '{default: 0};
        end
        else begin
            memory <= memory_next;
        end
    end

    parameter WORD_PER_BULK = 2**(WORD_ADDR_WIDTH-BULK_ADDR_WIDTH);

    logic [AGU_BITWIDTH-1:0] stages;
    logic [AGU_BITWIDTH-1:0] n_points;

    int i;
    always_comb begin
        if (fft_valid) begin
            n_points = n_points_0_0;
            stages = '0;
            for (i = AGU_BITWIDTH-1; i >= 0; i--) begin
                if (n_points[i]) begin
                    stages = i;
                    break;
                end
            end
        end
    end
    
    logic [WORD_ADDR_WIDTH-BULK_ADDR_WIDTH-1:0] offset_w_addr, offset_r_addr;

    // LUT with bit reversed sequence for bulk address read
    typedef bit [AGU_BITWIDTH-1:0] LUT_t [RF_DEPTH];

    function LUT_t LUT_init();
        LUT_t temp;
        logic [AGU_BITWIDTH*2-1:0] ref_addr;
        int j;
        
        foreach (temp[i]) begin
            ref_addr = i << AGU_BITWIDTH;
            // Bit reversal
            for (j = 0; j < AGU_BITWIDTH; j++) begin
                temp[i][j] = ref_addr[stages - 1 - j + AGU_BITWIDTH];
            end
        end
        
        return temp;
    endfunction

    LUT_t bit_rev_addr;
    // initial bit_rev_addr = LUT_init();
    
    always_comb begin
        memory_next = memory;
        bulk_data_out_0 = 0;
        word_data_out_0 = 0;
        word_data_out_1 = 0;
        if (bulk_w_en) begin
            for (int i=0; i<WORD_PER_BULK; i++) begin
                offset_w_addr = i;
                memory_next[{bulk_w_addr, offset_w_addr}] = bulk_data_in_0[i*WORD_BITWIDTH +:WORD_BITWIDTH];
            end
        end
        if (word_w_en_0) begin
            if ((!bulk_w_en) || (bulk_w_addr != word_w_addr_0[WORD_ADDR_WIDTH-1:WORD_ADDR_WIDTH-1-BULK_ADDR_WIDTH]) || word_w_addr_1 != word_w_addr_0) begin
                memory_next[word_w_addr_0] = word_data_in_0;
            end
        end
        if (word_w_en_1) begin
            if ((!bulk_w_en) || (bulk_w_addr != word_w_addr_1[WORD_ADDR_WIDTH-1:WORD_ADDR_WIDTH-1-BULK_ADDR_WIDTH]) || word_w_addr_0!= word_w_addr_1) begin
                memory_next[word_w_addr_1] = word_data_in_1;
            end
        end
        if (bulk_r_en) begin
            bit_rev_addr = LUT_init();
            for (int i=0; i<WORD_PER_BULK; i++) begin
                bulk_data_out_0[i*WORD_BITWIDTH +:WORD_BITWIDTH] = memory[bit_rev_addr[i+bulk_r_addr*WORD_PER_BULK]];
            end
        end
        if (word_r_en_0) begin
            word_data_out_0 = memory[word_r_addr_0];
        end
        if (word_r_en_1) begin
            word_data_out_1 = memory[word_r_addr_1];
        end

    end

    logic [INSTR_OPCODE_BITWIDTH-1:0] opcode;
    logic [RESOURCE_INSTR_WIDTH-INSTR_OPCODE_BITWIDTH-1:0] payload;

    assign opcode = instr_0[RESOURCE_INSTR_WIDTH-1:RESOURCE_INSTR_WIDTH-INSTR_OPCODE_BITWIDTH];
    assign payload = instr_0[RESOURCE_INSTR_WIDTH-INSTR_OPCODE_BITWIDTH-1:0];

    fft_t fft;
    dsu_t dsu;
    rep_t rep;

    assign dsu_valid = instr_en_0 && (opcode == 6);
    assign rep_valid = instr_en_0 && (opcode == 0);
    assign fft_valid = instr_en_0 && (opcode == 4);
    assign dsu = dsu_valid ? unpack_dsu(payload) : '{default: 0};
    assign rep = rep_valid ? unpack_rep(payload) : '{default: 0};
    assign fft = fft_valid ? unpack_fft(payload) : '{default: 0};

    assign n_points_0_0 = fft._n_points;
    assign radix_0_0 = fft._radix;
    assign mode_0_0 = fft._mode;
    assign n_bu_0_0 = fft._n_bu;
    assign delay_0_0 = fft._delay;
    assign n_points_0_1 = fft._n_points;
    assign radix_0_1 = fft._radix;
    assign mode_0_1 = fft._mode;
    assign n_bu_0_1 = fft._n_bu;
    assign delay_0_1 = fft._delay;

    assign step_0_2 = rep._step;
    assign delay_0_2 = rep._delay;
    assign iter_0_2 = rep._iter;
    assign init_addr_0_2 = dsu._init_addr;
    assign step_0_3 = rep._step;
    assign delay_0_3 = rep._delay;
    assign iter_0_3 = rep._iter;
    assign init_addr_0_3 = dsu._init_addr;

    assign n_points_1_0 = fft._n_points;
    assign radix_1_0 = fft._radix;
    assign mode_1_0 = fft._mode;
    assign n_bu_1_0 = fft._n_bu;
    assign delay_1_0 = fft._delay;
    assign n_points_1_1 = fft._n_points;
    assign radix_1_1 = fft._radix;
    assign mode_1_1 = fft._mode;
    assign n_bu_1_1 = fft._n_bu;
    assign delay_1_1 = fft._delay;

    agu_fft4 #(
        .AGU_BITWIDTH(AGU_BITWIDTH),
        .DELAY_WIDTH(DELAY_WIDTH)
    ) agu_0_0 (
        .clk(clk),
        .rst_n(rst_n),
        .activate(activate_0[0]),
        .radix(radix_0_0),
        .even_odd(1'b0),
        .mode(mode_0_0),
        .n_bu(n_bu_0_0),
        .bu_index(1'b0),
        .n_points(n_points_0_0),
        .delay(delay_0_0),
        .load_config(fft_valid & fft._port == 0),
        .address_valid(word_w_en_0),
        .address(word_w_agu_0)
    );

    agu_fft4 #(
        .AGU_BITWIDTH(AGU_BITWIDTH),
        .DELAY_WIDTH(DELAY_WIDTH)
    ) agu_0_1 (
        .clk(clk),
        .rst_n(rst_n),
        .activate(activate_0[1]),
        .radix(radix_0_1),
        .even_odd(1'b0),
        .mode(mode_0_1),
        .n_bu(n_bu_0_1),
        .bu_index(1'b0),
        .n_points(n_points_0_1),
        .delay(delay_0_1),
        .load_config(fft_valid & fft._port == 1),
        .address_valid(word_r_en_0),
        .address(word_r_agu_0)
    );

    agu #(
        .ADDRESS_WIDTH(AGU_BITWIDTH),
        .NUMBER_OF_LEVELS(4)
    ) agu_0_2 (
        .clk(clk),
        .rst_n(rst_n),
        .activate(activate_0[2]),
        .load_initial(dsu_valid & dsu._port == 2),
        .load_level(rep_valid & rep._port == 2),
        .is_extended(),  // TODO: not supported yet
        .level_to_load(rep._level[1:0]),
        .step(step_0_2),
        .delay(delay_0_2),
        .iterations(iter_0_2),
        .initial_address(init_addr_0_2),
        .address_valid(bulk_w_en),
        .address(bulk_w_agu)
    );

    agu #(
        .ADDRESS_WIDTH(AGU_BITWIDTH),
        .NUMBER_OF_LEVELS(4)
    ) agu_0_3 (
        .clk(clk),
        .rst_n(rst_n),
        .activate(activate_0[3]),
        .load_initial(dsu_valid & dsu._port == 3),
        .load_level(rep_valid & rep._port == 3),
        .is_extended(),  // TODO: not supported yet
        .level_to_load(rep._level[1:0]),
        .step(step_0_3),
        .delay(delay_0_3),
        .iterations(iter_0_3),
        .initial_address(init_addr_0_3),
        .address_valid(bulk_r_en),
        .address(bulk_r_agu)
    );

    agu_fft4 #(
        .AGU_BITWIDTH(AGU_BITWIDTH),
        .DELAY_WIDTH(DELAY_WIDTH)
    ) agu_1_0 (
        .clk(clk),
        .rst_n(rst_n),
        .activate(activate_1[0]),
        .radix(radix_1_0),
        .even_odd(1'b1),
        .mode(mode_1_0),
        .n_bu(n_bu_1_0),
        .bu_index(1'b1),
        .n_points(n_points_1_0),
        .delay(delay_1_0),
        .load_config(fft_valid & fft._port == 0),
        .address_valid(word_w_en_1),
        .address(word_w_agu_1)
    );

    agu_fft4 #(
        .AGU_BITWIDTH(AGU_BITWIDTH),
        .DELAY_WIDTH(DELAY_WIDTH)
    ) agu_1_1 (
        .clk(clk),
        .rst_n(rst_n),
        .activate(activate_1[1]),
        .radix(radix_1_1),
        .even_odd(1'b1),
        .mode(mode_1_1),
        .n_bu(n_bu_1_1),
        .bu_index(1'b1),
        .n_points(n_points_1_1),
        .delay(delay_1_1),
        .load_config(fft_valid & fft._port == 1),
        .address_valid(word_r_en_1),
        .address(word_r_agu_1)
    );

endmodule

