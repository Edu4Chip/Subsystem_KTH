`define cell_btm_impl _3cb39fcneue
`define cell_btm_impl_pkg _3cb39fcneue_pkg
`define cell_mid_impl _teewgpcaalx
`define cell_mid_impl_pkg _teewgpcaalx_pkg
`define cell_top_impl _gh3m7x647ap
`define cell_top_impl_pkg _gh3m7x647ap_pkg
`define complex_dpu_impl _uvcilbfxawa
`define complex_dpu_impl_pkg _uvcilbfxawa_pkg
`define iosram_btm_impl _hez9qsj1kug
`define iosram_btm_impl_pkg _hez9qsj1kug_pkg
`define iosram_top_impl _xbvdm4fjuts
`define iosram_top_impl_pkg _xbvdm4fjuts_pkg
`define radix2_bu_impl _geetgwgvwme
`define radix2_bu_impl_pkg _geetgwgvwme_pkg
`define rf_fft_impl _hxfcpuabvjh
`define rf_fft_impl_pkg _hxfcpuabvjh_pkg
`define sequencer_impl _bofiw7zs7vj
`define sequencer_impl_pkg _bofiw7zs7vj_pkg
`define swb_impl _dixk93xtnmt
`define swb_impl_pkg _dixk93xtnmt_pkg

package fabric_pkg;
    parameter BULK_WIDTH = 256;
    parameter COLS = 1;
    parameter INSTR_ADDR_WIDTH = 6;
    parameter INSTR_DATA_WIDTH = 32;
    parameter INSTR_HOPS_WIDTH = 4;
    parameter INSTR_OPCODE_BITWIDTH = 3;
    parameter IO_ADDR_WIDTH = 16;
    parameter IO_DATA_WIDTH = 256;
    parameter RESOURCE_INSTR_WIDTH = 27;
    parameter ROWS = 3;
endpackage

module fabric
import fabric_pkg::*;
(
    input  logic clk,
    input  logic rst_n,
    input  logic [ROWS-1:0] call,
    output logic [ROWS-1:0] ret,
    output logic [COLS-1:0] io_en_in,
    output logic [COLS-1:0][IO_ADDR_WIDTH-1:0] io_addr_in,
    input  logic [COLS-1:0][IO_DATA_WIDTH-1:0] io_data_in,
    output logic [COLS-1:0] io_en_out,
    output logic [COLS-1:0][IO_ADDR_WIDTH-1:0] io_addr_out,
    output logic [COLS-1:0][IO_DATA_WIDTH-1:0] io_data_out,
    input  logic [ROWS-1:0][INSTR_DATA_WIDTH-1:0] instr_data_in,
    input  logic [ROWS-1:0][INSTR_ADDR_WIDTH-1:0] instr_addr_in,
    input  logic [ROWS-1:0][INSTR_HOPS_WIDTH-1:0] instr_hops_in,
    input  logic [ROWS-1:0] instr_en_in,
    output logic [ROWS-1:0][INSTR_DATA_WIDTH-1:0] instr_data_out,
    output logic [ROWS-1:0][INSTR_ADDR_WIDTH-1:0] instr_addr_out,
    output logic [ROWS-1:0][INSTR_HOPS_WIDTH-1:0] instr_hops_out,
    output logic [ROWS-1:0] instr_en_out
);

    logic [ROWS-1:0][COLS:0] call_net;
    logic [ROWS-1:0][COLS:0] ret_net;
    logic [ROWS-1:0][COLS:0][INSTR_DATA_WIDTH-1:0] instr_data_net;
    logic [ROWS-1:0][COLS:0][INSTR_ADDR_WIDTH-1:0] instr_addr_net;
    logic [ROWS-1:0][COLS:0][INSTR_HOPS_WIDTH-1:0] instr_hops_net;
    logic [ROWS-1:0][COLS:0] instr_en_net;

    logic[ROWS:0][COLS:0][BULK_WIDTH-1:0] bulk_intercell_n2s_net;
    logic[ROWS:0][COLS:0][BULK_WIDTH-1:0] bulk_intercell_w2e_net;
    logic[ROWS:0][COLS:0][BULK_WIDTH-1:0] bulk_intercell_s2n_net;
    logic[ROWS:0][COLS:0][BULK_WIDTH-1:0] bulk_intercell_e2w_net;

    for(genvar i=0; i<ROWS; i++) begin
        assign ret[i] = ret_net[i][0];
        assign ret_net[i][COLS] = 1;
        assign call_net[i][0] = call[i];
        assign instr_data_net[i][0] = instr_data_in[i];
        assign instr_addr_net[i][0] = instr_addr_in[i];
        assign instr_hops_net[i][0] = instr_hops_in[i];
        assign instr_en_net[i][0] = instr_en_in[i];
        assign instr_data_out[i] = instr_data_net[i][COLS];
        assign instr_addr_out[i] = instr_addr_net[i][COLS];
        assign instr_hops_out[i] = instr_hops_net[i][COLS];
        assign instr_en_out[i] = instr_en_net[i][COLS];
    end
`cell_top_impl cell_0_0_inst (
        .clk(clk),
        .rst_n(rst_n),
        .call_in(call_net[0][0]),
        .call_out(call_net[0][1]),
        .ret_in(ret_net[0][1]),
        .ret_out(ret_net[0][0]),
        .io_en_in(io_en_in[0]),
        .io_addr_in(io_addr_in[0]),
        .io_data_in(io_data_in[0]),
        .instr_data_in(instr_data_net[0][0]),
        .instr_addr_in(instr_addr_net[0][0]),
        .instr_hops_in(instr_hops_net[0][0]),
        .instr_en_in(instr_en_net[0][0]),
        .instr_data_out(instr_data_net[0][1]),
        .instr_addr_out(instr_addr_net[0][1]),
        .instr_hops_out(instr_hops_net[0][1]),
        .instr_en_out(instr_en_net[0][1]),
        .bulk_intercell_n_in(bulk_intercell_n2s_net[0][0]),
        .bulk_intercell_w_in(bulk_intercell_w2e_net[0][0]),
        .bulk_intercell_s_in(bulk_intercell_s2n_net[1][0]),
        .bulk_intercell_e_in(bulk_intercell_e2w_net[0][1]),
        .bulk_intercell_n_out(bulk_intercell_s2n_net[0][0]),
        .bulk_intercell_w_out(bulk_intercell_w2e_net[0][0]),
        .bulk_intercell_s_out(bulk_intercell_n2s_net[1][0]),
        .bulk_intercell_e_out(bulk_intercell_e2w_net[0][1])
    );
`cell_mid_impl cell_1_0_inst (
        .clk(clk),
        .rst_n(rst_n),
        .call_in(call_net[1][0]),
        .call_out(call_net[1][1]),
        .ret_in(ret_net[1][1]),
        .ret_out(ret_net[1][0]),
        .io_data_in(io_data_in[0]),
        .instr_data_in(instr_data_net[1][0]),
        .instr_addr_in(instr_addr_net[1][0]),
        .instr_hops_in(instr_hops_net[1][0]),
        .instr_en_in(instr_en_net[1][0]),
        .instr_data_out(instr_data_net[1][1]),
        .instr_addr_out(instr_addr_net[1][1]),
        .instr_hops_out(instr_hops_net[1][1]),
        .instr_en_out(instr_en_net[1][1]),
        .bulk_intercell_n_in(bulk_intercell_n2s_net[1][0]),
        .bulk_intercell_w_in(bulk_intercell_w2e_net[1][0]),
        .bulk_intercell_s_in(bulk_intercell_s2n_net[2][0]),
        .bulk_intercell_e_in(bulk_intercell_e2w_net[1][1]),
        .bulk_intercell_n_out(bulk_intercell_s2n_net[1][0]),
        .bulk_intercell_w_out(bulk_intercell_w2e_net[1][0]),
        .bulk_intercell_s_out(bulk_intercell_n2s_net[2][0]),
        .bulk_intercell_e_out(bulk_intercell_e2w_net[1][1])
    );
`cell_btm_impl cell_2_0_inst (
        .clk(clk),
        .rst_n(rst_n),
        .call_in(call_net[2][0]),
        .call_out(call_net[2][1]),
        .ret_in(ret_net[2][1]),
        .ret_out(ret_net[2][0]),
        .io_data_in(io_data_in[0]),
        .io_en_out(io_en_out[0]),
        .io_addr_out(io_addr_out[0]),
        .io_data_out(io_data_out[0]),
        .instr_data_in(instr_data_net[2][0]),
        .instr_addr_in(instr_addr_net[2][0]),
        .instr_hops_in(instr_hops_net[2][0]),
        .instr_en_in(instr_en_net[2][0]),
        .instr_data_out(instr_data_net[2][1]),
        .instr_addr_out(instr_addr_net[2][1]),
        .instr_hops_out(instr_hops_net[2][1]),
        .instr_en_out(instr_en_net[2][1]),
        .bulk_intercell_n_in(bulk_intercell_n2s_net[2][0]),
        .bulk_intercell_w_in(bulk_intercell_w2e_net[2][0]),
        .bulk_intercell_s_in(bulk_intercell_s2n_net[3][0]),
        .bulk_intercell_e_in(bulk_intercell_e2w_net[2][1]),
        .bulk_intercell_n_out(bulk_intercell_s2n_net[2][0]),
        .bulk_intercell_w_out(bulk_intercell_w2e_net[2][0]),
        .bulk_intercell_s_out(bulk_intercell_n2s_net[3][0]),
        .bulk_intercell_e_out(bulk_intercell_e2w_net[2][1])
    );
endmodule