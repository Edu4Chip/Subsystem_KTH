`define sequencer_impl _bofiw7zs7vj
`define sequencer_impl_pkg _bofiw7zs7vj_pkg

package _bofiw7zs7vj_pkg;
    parameter FSM_PER_SLOT = 4;
    parameter INSTR_ADDR_WIDTH = 6;
    parameter INSTR_DATA_WIDTH = 32;
    parameter INSTR_HOPS_WIDTH = 4;
    parameter NUM_SLOTS = 16;
    parameter RESOURCE_INSTR_WIDTH = 27;

    // Others:
    typedef struct packed {
        logic _mode;
        logic [26:0] _cycle;
    } wait_t;

    function static wait_t unpack_wait;
        input logic [27:0] instr;
        wait_t _wait;
        _wait._mode = instr[27];
        _wait._cycle  = instr[26:0];
        return _wait;
    endfunction

    function static logic [27:0] pack_wait;
        input wait_t _wait;
        logic [27:0] instr;

        instr[27] = _wait._mode;
        instr[26:0] = _wait._cycle;
        return instr;
    endfunction
    typedef struct packed {
        logic [15:0] _ports;
        logic [3:0] _mode;
        logic [7:0] _param;
    } act_t;

    function static act_t unpack_act;
        input logic [27:0] instr;
        act_t _act;
        _act._ports  = instr[27:12];
        _act._mode  = instr[11:8];
        _act._param  = instr[7:0];
        return _act;
    endfunction

    function static logic [27:0] pack_act;
        input act_t _act;
        logic [27:0] instr;

        instr[27:12] = _act._ports;
        instr[11:8] = _act._mode;
        instr[7:0] = _act._param;
        return instr;
    endfunction
    typedef struct packed {
        logic [5:0] _mode;
        logic [3:0] _operand1;
        logic _operand2_sd;
        logic [7:0] _operand2;
        logic [3:0] _result;
    } calc_t;

    function static calc_t unpack_calc;
        input logic [27:0] instr;
        calc_t _calc;
        _calc._mode  = instr[27:22];
        _calc._operand1  = instr[21:18];
        _calc._operand2_sd = instr[17];
        _calc._operand2  = instr[16:9];
        _calc._result  = instr[8:5];
        return _calc;
    endfunction

    function static logic [27:0] pack_calc;
        input calc_t _calc;
        logic [27:0] instr;

        instr[27:22] = _calc._mode;
        instr[21:18] = _calc._operand1;
        instr[17] = _calc._operand2_sd;
        instr[16:9] = _calc._operand2;
        instr[8:5] = _calc._result;
        return instr;
    endfunction
    typedef struct packed {
        logic [3:0] _reg;
        logic [8:0] _target_true;
        logic [8:0] _target_false;
    } brn_t;

    function static brn_t unpack_brn;
        input logic [27:0] instr;
        brn_t _brn;
        _brn._reg  = instr[27:24];
        _brn._target_true  = instr[23:15];
        _brn._target_false  = instr[14:6];
        return _brn;
    endfunction

    function static logic [27:0] pack_brn;
        input brn_t _brn;
        logic [27:0] instr;

        instr[27:24] = _brn._reg;
        instr[23:15] = _brn._target_true;
        instr[14:6] = _brn._target_false;
        return instr;
    endfunction

endpackage
module _bofiw7zs7vj
import _bofiw7zs7vj_pkg::*;
(
    input  logic clk,
    input  logic rst_n,
    input  logic call,
    output logic ret,
    output logic instr_valid_0,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_0,
    output logic [FSM_PER_SLOT-1:0] activate_0,
    output logic clk_0,
    output logic rst_n_0,
    output logic instr_valid_1,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_1,
    output logic [FSM_PER_SLOT-1:0] activate_1,
    output logic clk_1,
    output logic rst_n_1,
    output logic instr_valid_2,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_2,
    output logic [FSM_PER_SLOT-1:0] activate_2,
    output logic clk_2,
    output logic rst_n_2,
    output logic instr_valid_3,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_3,
    output logic [FSM_PER_SLOT-1:0] activate_3,
    output logic clk_3,
    output logic rst_n_3,
    output logic instr_valid_4,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_4,
    output logic [FSM_PER_SLOT-1:0] activate_4,
    output logic clk_4,
    output logic rst_n_4,
    output logic instr_valid_5,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_5,
    output logic [FSM_PER_SLOT-1:0] activate_5,
    output logic clk_5,
    output logic rst_n_5,
    output logic instr_valid_6,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_6,
    output logic [FSM_PER_SLOT-1:0] activate_6,
    output logic clk_6,
    output logic rst_n_6,
    output logic instr_valid_7,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_7,
    output logic [FSM_PER_SLOT-1:0] activate_7,
    output logic clk_7,
    output logic rst_n_7,
    output logic instr_valid_8,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_8,
    output logic [FSM_PER_SLOT-1:0] activate_8,
    output logic clk_8,
    output logic rst_n_8,
    output logic instr_valid_9,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_9,
    output logic [FSM_PER_SLOT-1:0] activate_9,
    output logic clk_9,
    output logic rst_n_9,
    output logic instr_valid_10,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_10,
    output logic [FSM_PER_SLOT-1:0] activate_10,
    output logic clk_10,
    output logic rst_n_10,
    output logic instr_valid_11,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_11,
    output logic [FSM_PER_SLOT-1:0] activate_11,
    output logic clk_11,
    output logic rst_n_11,
    output logic instr_valid_12,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_12,
    output logic [FSM_PER_SLOT-1:0] activate_12,
    output logic clk_12,
    output logic rst_n_12,
    output logic instr_valid_13,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_13,
    output logic [FSM_PER_SLOT-1:0] activate_13,
    output logic clk_13,
    output logic rst_n_13,
    output logic instr_valid_14,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_14,
    output logic [FSM_PER_SLOT-1:0] activate_14,
    output logic clk_14,
    output logic rst_n_14,
    output logic instr_valid_15,
    output logic [RESOURCE_INSTR_WIDTH-1:0] instr_15,
    output logic [FSM_PER_SLOT-1:0] activate_15,
    output logic clk_15,
    output logic rst_n_15,
    input  logic [INSTR_DATA_WIDTH-1:0] instr_load_data_in,
    input  logic [INSTR_ADDR_WIDTH-1:0] instr_load_addr_in,
    input  logic [INSTR_HOPS_WIDTH-1:0] instr_load_hops_in,
    input  logic instr_load_en_in,
    output logic [INSTR_DATA_WIDTH-1:0] instr_load_data_out,
    output logic [INSTR_ADDR_WIDTH-1:0] instr_load_addr_out,
    output logic [INSTR_HOPS_WIDTH-1:0] instr_load_hops_out,
    output logic instr_load_en_out
);

    // Propagate signals to resources:
    logic [NUM_SLOTS-1:0] resource_instr;
    logic [RESOURCE_INSTR_WIDTH-1:0] instr;
    logic [NUM_SLOTS-1:0] resource_instr_valid;
    logic [NUM_SLOTS-1:0][FSM_PER_SLOT-1:0] resource_activate;
    assign clk_0 = clk;
    assign rst_n_0 = rst_n;
    assign instr_valid_0 = resource_instr_valid[0];
    assign activate_0 = resource_activate[0];
    assign instr_0 = instr;
    assign clk_1 = clk;
    assign rst_n_1 = rst_n;
    assign instr_valid_1 = resource_instr_valid[1];
    assign activate_1 = resource_activate[1];
    assign instr_1 = instr;
    assign clk_2 = clk;
    assign rst_n_2 = rst_n;
    assign instr_valid_2 = resource_instr_valid[2];
    assign activate_2 = resource_activate[2];
    assign instr_2 = instr;
    assign clk_3 = clk;
    assign rst_n_3 = rst_n;
    assign instr_valid_3 = resource_instr_valid[3];
    assign activate_3 = resource_activate[3];
    assign instr_3 = instr;
    assign clk_4 = clk;
    assign rst_n_4 = rst_n;
    assign instr_valid_4 = resource_instr_valid[4];
    assign activate_4 = resource_activate[4];
    assign instr_4 = instr;
    assign clk_5 = clk;
    assign rst_n_5 = rst_n;
    assign instr_valid_5 = resource_instr_valid[5];
    assign activate_5 = resource_activate[5];
    assign instr_5 = instr;
    assign clk_6 = clk;
    assign rst_n_6 = rst_n;
    assign instr_valid_6 = resource_instr_valid[6];
    assign activate_6 = resource_activate[6];
    assign instr_6 = instr;
    assign clk_7 = clk;
    assign rst_n_7 = rst_n;
    assign instr_valid_7 = resource_instr_valid[7];
    assign activate_7 = resource_activate[7];
    assign instr_7 = instr;
    assign clk_8 = clk;
    assign rst_n_8 = rst_n;
    assign instr_valid_8 = resource_instr_valid[8];
    assign activate_8 = resource_activate[8];
    assign instr_8 = instr;
    assign clk_9 = clk;
    assign rst_n_9 = rst_n;
    assign instr_valid_9 = resource_instr_valid[9];
    assign activate_9 = resource_activate[9];
    assign instr_9 = instr;
    assign clk_10 = clk;
    assign rst_n_10 = rst_n;
    assign instr_valid_10 = resource_instr_valid[10];
    assign activate_10 = resource_activate[10];
    assign instr_10 = instr;
    assign clk_11 = clk;
    assign rst_n_11 = rst_n;
    assign instr_valid_11 = resource_instr_valid[11];
    assign activate_11 = resource_activate[11];
    assign instr_11 = instr;
    assign clk_12 = clk;
    assign rst_n_12 = rst_n;
    assign instr_valid_12 = resource_instr_valid[12];
    assign activate_12 = resource_activate[12];
    assign instr_12 = instr;
    assign clk_13 = clk;
    assign rst_n_13 = rst_n;
    assign instr_valid_13 = resource_instr_valid[13];
    assign activate_13 = resource_activate[13];
    assign instr_13 = instr;
    assign clk_14 = clk;
    assign rst_n_14 = rst_n;
    assign instr_valid_14 = resource_instr_valid[14];
    assign activate_14 = resource_activate[14];
    assign instr_14 = instr;
    assign clk_15 = clk;
    assign rst_n_15 = rst_n;
    assign instr_valid_15 = resource_instr_valid[15];
    assign activate_15 = resource_activate[15];
    assign instr_15 = instr;

    // Parameter check:

    // Function definition:
    logic [NUM_SLOTS * FSM_PER_SLOT - 1:0] activate_flat;

    logic [27:0] instr_reg;
    logic [63:0][31:0] iram;
    logic [3:0] opcode;
    logic instr_type;
    logic [3:0] slot;
    logic [23:0] payload;
    logic [5:0] pc, pc_next;
    logic [16:0] wait_counter, wait_counter_next;

    typedef enum logic [1:0] { RESET, IDLE, DECODE, WAIT} state_t;
    state_t state, next_state;

    assign instr_type = iram[pc][31];
    assign opcode = iram[pc][30:28];
    assign instr_reg = iram[pc][27:0];
    assign payload = iram[pc][23:0];
    assign slot = iram[pc][27:24];

    always_ff @(posedge clk or negedge rst_n) begin
        if (~rst_n) begin
            instr_load_data_out <= 0;
            instr_load_addr_out <= 0;
            instr_load_hops_out <= 0;
            instr_load_en_out <= 0;
            for (int i=0; i<64; i++) begin
                iram[i] <= 0;
            end
        end else begin
            if (instr_load_en_in) begin
                if (instr_load_hops_in == 0) begin
                    iram[instr_load_addr_in] <= instr_load_data_in;
                    instr_load_data_out <= 0;
                    instr_load_addr_out <= 0;
                    instr_load_hops_out <= 0;
                    instr_load_en_out <= 0;
                end else begin
                    instr_load_data_out <= instr_load_data_in;
                    instr_load_addr_out <= instr_load_addr_in;
                    instr_load_hops_out <= instr_load_hops_in - 1;
                    instr_load_en_out <= instr_load_en_in;
                end
            end else begin
                instr_load_data_out <= 0;
                instr_load_addr_out <= 0;
                instr_load_hops_out <= 0;
                instr_load_en_out <= 0;
            end
        end
    end

    // FSM:
    always_ff @(posedge clk or negedge rst_n) begin
        if (~rst_n) begin
            state <= RESET;
            pc <= 0;
            wait_counter <= 0;
        end else begin
            state <= next_state;
            pc <= pc_next;
            wait_counter <= wait_counter_next;
        end
    end

    always_comb begin
        next_state = state;
        pc_next = pc+1;
        wait_counter_next = wait_counter;
        case (state)
            RESET: begin
                next_state = IDLE;
                pc_next = 0;
            end
            IDLE: begin
                if (call == 1) begin
                    next_state = DECODE;
                    pc_next = 0;
                end else begin
                    next_state = IDLE;
                    pc_next = 0;
                end
            end
            DECODE: begin
                if (instr_type == 0 && opcode == 0) begin
                    pc_next = 0;
                    next_state = IDLE;
                end else if (instr_type == 0 && opcode == 1) begin
                    wait_t _wait;
                    _wait = unpack_wait(instr_reg);
                    if (_wait._cycle != 0) begin
                        pc_next = pc;
                        next_state = WAIT;
                        wait_counter_next = _wait._cycle;
                    end
                end
            end
            WAIT: begin
                wait_counter_next = wait_counter - 1;
                if (wait_counter == 1) begin
                    next_state = DECODE;
                end else begin
                    next_state = WAIT;
                    pc_next = pc;
                end
            end
        endcase
    end

    act_t _act;
    always_comb begin
        ret = 0;
        for (int i = 0; i < NUM_SLOTS; i = i + 1) begin
            resource_instr_valid[i] = 0;
            resource_activate[i] = 0;
        end
        instr = 0;
        case (state)
            DECODE: begin
                if (instr_type == 0) begin
                    if (opcode == 2) begin
                        activate_flat = 0;
                        _act = unpack_act(instr_reg);
                        activate_flat = _act._ports << (_act._param * FSM_PER_SLOT);
                        for (int i=0; i<NUM_SLOTS; i++) begin
                            resource_activate[i] = activate_flat[FSM_PER_SLOT*i +: FSM_PER_SLOT];
                        end
                    end else if (opcode == 0) begin
                        ret = 1;
                    end
                end else begin
                    instr = {opcode, payload};
                    resource_instr_valid[slot] = 1;
                end
            end
        endcase
    end
endmodule

